-- megafunction wizard: %Serial Flash Loader%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altserial_flash_loader 

-- ============================================================
-- File Name: ADV_SFL.vhd
-- Megafunction Name(s):
-- 			altserial_flash_loader
--
-- Simulation Library Files(s):
-- 			altera_mf
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 13.1.4 Build 182 03/12/2014 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2014 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY altera_mf;
USE altera_mf.all;

ENTITY ADV_SFL IS
	PORT
	(
		asdo_in		: IN STD_LOGIC ;
		asmi_access_granted		: IN STD_LOGIC ;
		dclk_in		: IN STD_LOGIC ;
		ncso_in		: IN STD_LOGIC ;
		noe_in		: IN STD_LOGIC ;
		asmi_access_request		: OUT STD_LOGIC ;
		data0_out		: OUT STD_LOGIC 
	);
END ADV_SFL;


ARCHITECTURE SYN OF adv_sfl IS

	SIGNAL sub_wire0	: STD_LOGIC ;
	SIGNAL sub_wire1	: STD_LOGIC ;



	COMPONENT altserial_flash_loader
	GENERIC (
		enable_quad_spi_support		: NATURAL;
		enable_shared_access		: STRING;
		enhanced_mode		: NATURAL;
		intended_device_family		: STRING;
		lpm_type		: STRING
	);
	PORT (
			data0out	: OUT STD_LOGIC ;
			noe	: IN STD_LOGIC ;
			scein	: IN STD_LOGIC ;
			asmi_access_granted	: IN STD_LOGIC ;
			asmi_access_request	: OUT STD_LOGIC ;
			dclkin	: IN STD_LOGIC ;
			sdoin	: IN STD_LOGIC 
	);
	END COMPONENT;

BEGIN
	asmi_access_request    <= sub_wire0;
	data0_out    <= sub_wire1;

	altserial_flash_loader_component : altserial_flash_loader
	GENERIC MAP (
		enable_quad_spi_support => 0,
		enable_shared_access => "ON",
		enhanced_mode => 1,
		intended_device_family => "Cyclone IV GX",
		lpm_type => "altserial_flash_loader"
	)
	PORT MAP (
		noe => noe_in,
		scein => ncso_in,
		asmi_access_granted => asmi_access_granted,
		dclkin => dclk_in,
		sdoin => asdo_in,
		asmi_access_request => sub_wire0,
		data0out => sub_wire1
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV GX"
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: ENABLE_QUAD_SPI_SUPPORT NUMERIC "0"
-- Retrieval info: CONSTANT: ENABLE_SHARED_ACCESS STRING "ON"
-- Retrieval info: CONSTANT: ENHANCED_MODE NUMERIC "1"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone IV GX"
-- Retrieval info: USED_PORT: asdo_in 0 0 0 0 INPUT NODEFVAL "asdo_in"
-- Retrieval info: USED_PORT: asmi_access_granted 0 0 0 0 INPUT NODEFVAL "asmi_access_granted"
-- Retrieval info: USED_PORT: asmi_access_request 0 0 0 0 OUTPUT NODEFVAL "asmi_access_request"
-- Retrieval info: USED_PORT: data0_out 0 0 0 0 OUTPUT NODEFVAL "data0_out"
-- Retrieval info: USED_PORT: dclk_in 0 0 0 0 INPUT NODEFVAL "dclk_in"
-- Retrieval info: USED_PORT: ncso_in 0 0 0 0 INPUT NODEFVAL "ncso_in"
-- Retrieval info: USED_PORT: noe_in 0 0 0 0 INPUT NODEFVAL "noe_in"
-- Retrieval info: CONNECT: @asmi_access_granted 0 0 0 0 asmi_access_granted 0 0 0 0
-- Retrieval info: CONNECT: @dclkin 0 0 0 0 dclk_in 0 0 0 0
-- Retrieval info: CONNECT: @noe 0 0 0 0 noe_in 0 0 0 0
-- Retrieval info: CONNECT: @scein 0 0 0 0 ncso_in 0 0 0 0
-- Retrieval info: CONNECT: @sdoin 0 0 0 0 asdo_in 0 0 0 0
-- Retrieval info: CONNECT: asmi_access_request 0 0 0 0 @asmi_access_request 0 0 0 0
-- Retrieval info: CONNECT: data0_out 0 0 0 0 @data0out 0 0 0 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL ADV_SFL.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ADV_SFL.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ADV_SFL.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ADV_SFL.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ADV_SFL_inst.vhd FALSE
-- Retrieval info: LIB_FILE: altera_mf
